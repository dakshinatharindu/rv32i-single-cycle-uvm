package core_pkg;

    // uvm
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // uvm_object

    // uvm_transactions

    // uvm_subscribers

    // uvm_agents

    // uvm_environment

    // uvm_tests
    
endpackage